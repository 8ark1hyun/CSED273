/* CSED273 lab4 experiment 3 */
/* lab4_3.v */
/* 20220100 박기현 */

/* Implement 5-Bit Ripple Subtractor
 * You must use lab4_2 module in lab4_2.v
 * You may use keword "assign" and bitwise operator
 * or just implement with gate-level modeling*/
module lab4_3(
    input [4:0] in_a,
    input [4:0] in_b,
    input in_c,
    output [4:0] out_s,
    output out_c
    );

    ////////////////////////
    lab4_2 Adder (in_a, ~in_b, in_c, out_s, out_c);
    ////////////////////////

endmodule
/* CSED273 lab1 experiment 2_iii */
/* lab1_2_iii.v */
/* 20220100 박기현 */

module lab1_2_iii(outAND, outOR, outNOT, inA, inB);
    output wire outAND, outOR, outNOT;
    input wire inA, inB;

    AND(outAND, inA, inB);
    OR(outOR, inA, inB);
    NOT(outNOT, inA);

endmodule


/* Implement AND, OR, and NOT modules with {NAND}
 * You are only allowed to wire modules below
 * i.e.) No and, or, not, etc. Only nand, AND, OR, NOT are available*/
module AND(outAND, inA, inB);
    output wire outAND;
    input wire inA, inB; 

    ////////////////////////
    wire C;
    nand(C, inA, inB); //C = NOT(A AND B)
    nand(outAND, C, C); //A AND B
    ////////////////////////

endmodule

module OR(outOR, inA, inB);
    output wire outOR;
    input wire inA, inB; 
    
    ////////////////////////
    wire D, E;
    nand(D, inA, inA); //D = NOT A
    nand(E, inB, inB); //E = NOT B
    nand(outOR, D, E); //A OR B
    ////////////////////////

endmodule

module NOT(outNOT, inA);
    output wire outNOT;
    input wire inA; 

    ////////////////////////
    nand(outNOT, inA, inA); //NOT A
    ////////////////////////

endmodule